`include "alu.v"
module top (
    ports
);
    
endmodule

module dmem (
    input clk, input [31:0] MemWrite, input [31:0] ALUResult, [31:0] WriteData,
    output [31:0] ReadData
);
    
endmodule

module imem (
    ports
);
    
endmodule

module controller (
    ports
);
    
endmodule

module datapath (
    ports
);
    
endmodule

module decode (
    ports
);
    
endmodule

module condlogic (
    output RegWrite, MemWrite, PCSrc
);
    
endmodule

